`ifndef FPU_PKG_INC_SV
`define FPU_PKG_INC_SV

`include "data_type_pkg.sv"
`include "op_intf.sv"

`endif
