`ifndef FPU_PKG_INC_SVH
`define FPU_PKG_INC_SVH

`define MODE_WIDTH 4
`define DATA_WIDTH 16

`define MODE_ADD 4'b0001
`define MODE_SUB 4'b0010
`define MODE_MUL 4'b0100
`define MODE_DIV 4'b1000

`endif